module TAADDA (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(8'd0), .en(wire_53[0:0]), .out(arch_output_value));
  TC_Counter # (.UUID(64'd188627541998958090 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_1 (.clk(clk), .rst(rst), .save(wire_16[0:0]), .in(wire_32), .out(wire_43));
  TC_Splitter8 # (.UUID(64'd3798056121934110910 ^ UUID)) Splitter8_2 (.in(wire_44[7:0]), .out0(wire_59), .out1(wire_36), .out2(wire_78), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2763155547170517442 ^ UUID)) Decoder3_3 (.dis(1'd0), .sel0(wire_59), .sel1(wire_36), .sel2(wire_78), .out0(wire_79), .out1(wire_54), .out2(wire_33), .out3(wire_83), .out4(wire_60), .out5(wire_71), .out6(wire_29), .out7(wire_68));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_4 (.en(wire_76), .in(arch_input_value), .out(wire_51));
  TC_Splitter8 # (.UUID(64'd1378806238108263558 ^ UUID)) Splitter8_5 (.in(wire_58[7:0]), .out0(wire_7), .out1(wire_9), .out2(wire_73), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2132310256929947462 ^ UUID)) Decoder3_6 (.dis(1'd0), .sel0(wire_7), .sel1(wire_9), .sel2(wire_73), .out0(wire_26), .out1(wire_52), .out2(wire_82), .out3(wire_61), .out4(wire_47), .out5(wire_2), .out6(wire_6), .out7(wire_80));
  TC_Decoder3 # (.UUID(64'd1568863074849052991 ^ UUID)) Decoder3_7 (.dis(1'd0), .sel0(wire_21), .sel1(wire_77), .sel2(wire_48), .out0(wire_11), .out1(wire_64), .out2(wire_22), .out3(wire_28), .out4(wire_35), .out5(wire_49), .out6(wire_39), .out7(wire_74));
  TC_Splitter8 # (.UUID(64'd4565437463060912785 ^ UUID)) Splitter8_8 (.in(wire_65[7:0]), .out0(wire_21), .out1(wire_77), .out2(wire_48), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Constant # (.UUID(64'd664116279942053836 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out(wire_76));
  TC_Switch # (.UUID(64'd2622295034880516622 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_24[0:0]), .in(wire_51), .out(wire_40_6));
  TC_Switch # (.UUID(64'd268561600865225889 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_38[0:0]), .in(wire_51), .out(wire_12_7));
  TC_Switch # (.UUID(64'd2366302977062530316 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_13[0:0]), .in(wire_62), .out(wire_12_1));
  TC_Switch # (.UUID(64'd1161835394234352669 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_66[0:0]), .in(wire_62), .out(wire_40_5));
  TC_Switch # (.UUID(64'd664368396214293951 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_10[0:0]), .in(wire_45), .out(wire_12_0));
  TC_Switch # (.UUID(64'd971706953703219603 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_0[0:0]), .in(wire_45), .out(wire_40_3));
  TC_Switch # (.UUID(64'd550582960029639035 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_1[0:0]), .in(wire_27), .out(wire_12_2));
  TC_Switch # (.UUID(64'd2551371438056267438 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_17[0:0]), .in(wire_27), .out(wire_40_1));
  TC_Switch # (.UUID(64'd1328714823458733387 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_41[0:0]), .in(wire_63), .out(wire_12_3));
  TC_Switch # (.UUID(64'd4275065018319978774 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_50[0:0]), .in(wire_63), .out(wire_40_0));
  TC_Switch # (.UUID(64'd2071649843942799398 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_19[0:0]), .in(wire_5), .out(wire_12_5));
  TC_Switch # (.UUID(64'd1204434183799054386 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_69[0:0]), .in(wire_5), .out(wire_40_2));
  TC_Switch # (.UUID(64'd469546117461052876 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_42[0:0]), .in(wire_67), .out(wire_12_6));
  TC_Switch # (.UUID(64'd3273196033402958089 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_55[0:0]), .in(wire_67), .out(wire_40_4));
  TC_Switch # (.UUID(64'd3539769237345777454 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_23[0:0]), .in(wire_43), .out(wire_40_8));
  TC_Switch # (.UUID(64'd559995122624790222 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_31[0:0]), .in(wire_43), .out(wire_12_8));
  TC_Splitter8 # (.UUID(64'd3402866529736890305 ^ UUID)) Splitter8_26 (.in(wire_25[7:0]), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(wire_20), .out6(wire_57), .out7(wire_4));
  TC_Switch # (.UUID(64'd3278352177646989803 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_4), .in(wire_58[7:0]), .out(wire_12_4));
  TC_Switch # (.UUID(64'd2895273590468657512 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_57), .in(wire_65[7:0]), .out(wire_40_7));
  TC_Not # (.UUID(64'd2892521605633732722 ^ UUID), .BIT_WIDTH(64'd1)) Not_29 (.in(wire_57), .out(wire_14));
  TC_Not # (.UUID(64'd1891312441340278586 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_4), .out(wire_3));
  TC_Switch # (.UUID(64'd1244685540260459335 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_14), .in({{7{1'b0}}, wire_11 }), .out(wire_66));
  TC_Switch # (.UUID(64'd1077755302843490829 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_14), .in({{7{1'b0}}, wire_64 }), .out(wire_0));
  TC_Switch # (.UUID(64'd2165702842962589731 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_14), .in({{7{1'b0}}, wire_22 }), .out(wire_17));
  TC_Switch # (.UUID(64'd3617536616208170204 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_14), .in({{7{1'b0}}, wire_28 }), .out(wire_50));
  TC_Switch # (.UUID(64'd1296625335259484905 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_14), .in({{7{1'b0}}, wire_35 }), .out(wire_69));
  TC_Switch # (.UUID(64'd407289912901857071 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_14), .in({{7{1'b0}}, wire_49 }), .out(wire_55));
  TC_Switch # (.UUID(64'd3551958095488279259 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_37 (.en(wire_14), .in({{7{1'b0}}, wire_39 }), .out(wire_23));
  TC_Switch # (.UUID(64'd945374254991909364 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_14), .in({{7{1'b0}}, wire_74 }), .out(wire_24));
  TC_Switch # (.UUID(64'd2017577839392913570 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_39 (.en(wire_3), .in({{7{1'b0}}, wire_26 }), .out(wire_13));
  TC_Switch # (.UUID(64'd4222629416148848896 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_40 (.en(wire_3), .in({{7{1'b0}}, wire_52 }), .out(wire_10));
  TC_Switch # (.UUID(64'd956896318737315687 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_41 (.en(wire_3), .in({{7{1'b0}}, wire_82 }), .out(wire_1));
  TC_Switch # (.UUID(64'd2685356178464155659 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_3), .in({{7{1'b0}}, wire_61 }), .out(wire_41));
  TC_Switch # (.UUID(64'd2393103036448971650 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_3), .in({{7{1'b0}}, wire_47 }), .out(wire_19));
  TC_Switch # (.UUID(64'd2084091346705141896 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_3), .in({{7{1'b0}}, wire_2 }), .out(wire_42));
  TC_Switch # (.UUID(64'd4121630312737265200 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_3), .in({{7{1'b0}}, wire_6 }), .out(wire_31));
  TC_Switch # (.UUID(64'd4413701382283253951 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_3), .in({{7{1'b0}}, wire_80 }), .out(wire_38));
  TC_Switch # (.UUID(64'd3078506067986260760 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_15), .in({{7{1'b0}}, wire_79 }), .out(wire_75));
  TC_Switch # (.UUID(64'd4367250176294378390 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_15), .in({{7{1'b0}}, wire_54 }), .out(wire_56));
  TC_Switch # (.UUID(64'd125014847929148177 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_15), .in({{7{1'b0}}, wire_33 }), .out(wire_81));
  TC_Switch # (.UUID(64'd2927510286954144234 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_15), .in({{7{1'b0}}, wire_83 }), .out(wire_30));
  TC_Switch # (.UUID(64'd2252272992286407449 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_15), .in({{7{1'b0}}, wire_60 }), .out(wire_34));
  TC_Switch # (.UUID(64'd145110541831669376 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_15), .in({{7{1'b0}}, wire_71 }), .out(wire_8));
  TC_Switch # (.UUID(64'd3725212696777837935 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_15), .in({{7{1'b0}}, wire_29 }), .out(wire_16_1));
  TC_Switch # (.UUID(64'd4477946882270936064 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_15), .in({{7{1'b0}}, wire_68 }), .out(wire_53));
  TC_Not # (.UUID(64'd3879044616685914771 ^ UUID), .BIT_WIDTH(64'd1)) Not_55 (.in(wire_20), .out(wire_15));
  TC_Switch # (.UUID(64'd1942275899723426160 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_20), .in(wire_44[7:0]), .out(wire_46));
  TC_Switch # (.UUID(64'd1630534160172660904 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_37), .in(wire_46), .out(wire_32_0));
  TC_And # (.UUID(64'd1143668735634148691 ^ UUID), .BIT_WIDTH(64'd1)) And_58 (.in0(wire_18), .in1(wire_20), .out(wire_37));
  TC_Nand # (.UUID(64'd2856250237191538366 ^ UUID), .BIT_WIDTH(64'd1)) Nand_59 (.in0(wire_18), .in1(wire_20), .out(wire_72));
  TC_Switch # (.UUID(64'd865630561599775162 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_60 (.en(wire_72), .in({{7{1'b0}}, wire_18 }), .out(wire_32_1));
  TC_Switch # (.UUID(64'd2889242153891173726 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_61 (.en(wire_37), .in(wire_70), .out(wire_16_0[0:0]));
  TC_Constant # (.UUID(64'd2144963182158506193 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_62 (.out(wire_70));
  RegisterPlus # (.UUID(64'd4267416359963304908 ^ UUID)) RegisterPlus_63 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_8[0:0]), .Always_output(wire_67), .Output());
  RegisterPlus # (.UUID(64'd1069821230610740673 ^ UUID)) RegisterPlus_64 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_34[0:0]), .Always_output(wire_5), .Output());
  RegisterPlus # (.UUID(64'd1214749861541894319 ^ UUID)) RegisterPlus_65 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_30[0:0]), .Always_output(wire_63), .Output());
  RegisterPlus # (.UUID(64'd3854397592339658146 ^ UUID)) RegisterPlus_66 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_81[0:0]), .Always_output(wire_27), .Output());
  RegisterPlus # (.UUID(64'd773893054593625520 ^ UUID)) RegisterPlus_67 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_56[0:0]), .Always_output(wire_45), .Output());
  RegisterPlus # (.UUID(64'd4381960087344303846 ^ UUID)) RegisterPlus_68 (.clk(clk), .rst(rst), .Load(1'd0), .Save_value({{7{1'b0}}, wire_18 }), .Save(wire_75[0:0]), .Always_output(wire_62), .Output());
  TC_Program # (.UUID(64'd1175525504470668834 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_10504E37D662D622.w8.bin"), .ARG_SIG("Program_10504E37D662D622=%s")) Program_69 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_43 }), .out0(wire_25), .out1(wire_58), .out2(wire_65), .out3(wire_44));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_12_0;
  wire [7:0] wire_12_1;
  wire [7:0] wire_12_2;
  wire [7:0] wire_12_3;
  wire [7:0] wire_12_4;
  wire [7:0] wire_12_5;
  wire [7:0] wire_12_6;
  wire [7:0] wire_12_7;
  wire [7:0] wire_12_8;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2|wire_12_3|wire_12_4|wire_12_5|wire_12_6|wire_12_7|wire_12_8;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_16_0;
  wire [7:0] wire_16_1;
  assign wire_16 = wire_16_0|wire_16_1;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  assign wire_18 = 0;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_24;
  wire [63:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_32_0;
  wire [7:0] wire_32_1;
  assign wire_32 = wire_32_0|wire_32_1;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [7:0] wire_40_0;
  wire [7:0] wire_40_1;
  wire [7:0] wire_40_2;
  wire [7:0] wire_40_3;
  wire [7:0] wire_40_4;
  wire [7:0] wire_40_5;
  wire [7:0] wire_40_6;
  wire [7:0] wire_40_7;
  wire [7:0] wire_40_8;
  assign wire_40 = wire_40_0|wire_40_1|wire_40_2|wire_40_3|wire_40_4|wire_40_5|wire_40_6|wire_40_7|wire_40_8;
  wire [7:0] wire_41;
  wire [7:0] wire_42;
  wire [7:0] wire_43;
  wire [63:0] wire_44;
  wire [7:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [7:0] wire_53;
  assign arch_output_enable = wire_53[0:0];
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [0:0] wire_57;
  wire [63:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [7:0] wire_63;
  wire [0:0] wire_64;
  wire [63:0] wire_65;
  wire [7:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  assign arch_input_enable = wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;

endmodule
