module TAADDA (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_0), .en(wire_73), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_40), .in(arch_input_value), .out(wire_8));
  TC_Counter # (.UUID(64'd103235486555922174 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_2 (.clk(clk), .rst(rst), .save(wire_45), .in(wire_51), .out(wire_36));
  TC_Splitter8 # (.UUID(64'd278438544036793448 ^ UUID)) Splitter8_3 (.in(wire_86), .out0(wire_65), .out1(wire_87), .out2(wire_77), .out3(wire_6), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd1057399239572939361 ^ UUID)) Decoder3_4 (.dis(wire_17), .sel0(wire_65), .sel1(wire_87), .sel2(wire_77), .out0(wire_85), .out1(wire_82), .out2(wire_34), .out3(wire_49), .out4(wire_11), .out5(wire_29), .out6(wire_47), .out7(wire_73));
  TC_Splitter8 # (.UUID(64'd3708228715471769789 ^ UUID)) Splitter8_5 (.in(wire_5[7:0]), .out0(wire_80), .out1(wire_75), .out2(wire_83), .out3(wire_19), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd752126497560934249 ^ UUID)) Decoder3_6 (.dis(wire_19), .sel0(wire_80), .sel1(wire_75), .sel2(wire_83), .out0(wire_30), .out1(wire_84), .out2(wire_53), .out3(wire_37), .out4(wire_23), .out5(wire_24), .out6(wire_42), .out7(wire_39));
  TC_Decoder3 # (.UUID(64'd2653145962724689128 ^ UUID)) Decoder3_7 (.dis(wire_14), .sel0(wire_9), .sel1(wire_57), .sel2(wire_3), .out0(wire_81), .out1(wire_55), .out2(wire_67), .out3(wire_78), .out4(wire_26), .out5(wire_59), .out6(wire_20), .out7(wire_13));
  TC_Splitter8 # (.UUID(64'd2433189120953899482 ^ UUID)) Splitter8_8 (.in(wire_10[7:0]), .out0(wire_9), .out1(wire_57), .out2(wire_3), .out3(wire_14), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd1967783176326562294 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_13), .in(wire_8), .out(wire_4_7));
  TC_Switch # (.UUID(64'd1144500226581355342 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_39), .in(wire_8), .out(wire_28_1));
  TC_Switch # (.UUID(64'd4563522032870272540 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_42), .in(wire_36), .out(wire_28_7));
  TC_Switch # (.UUID(64'd1520248560007323449 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_20), .in(wire_36), .out(wire_4_2));
  TC_Mux # (.UUID(64'd4552121396603208012 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_13 (.sel(wire_16[0:0]), .in0(wire_4), .in1(wire_10[7:0]), .out(wire_58));
  TC_Mux # (.UUID(64'd1508906682506212572 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_14 (.sel(wire_18[0:0]), .in0(wire_28), .in1(wire_5[7:0]), .out(wire_1));
  TC_Splitter8 # (.UUID(64'd222548830488705950 ^ UUID)) Splitter8_15 (.in(wire_27[7:0]), .out0(wire_71), .out1(wire_60), .out2(wire_52), .out3(wire_22), .out4(), .out5(wire_35), .out6(), .out7());
  TC_Or # (.UUID(64'd3829124389360355821 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_47), .in1(wire_54), .out(wire_45));
  TC_Mux # (.UUID(64'd1711495082167809336 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_17 (.sel(wire_35), .in0(wire_0), .in1(wire_70), .out(wire_51));
  TC_And # (.UUID(64'd2465327194030448632 ^ UUID), .BIT_WIDTH(64'd1)) And_18 (.in0(wire_44), .in1(wire_35), .out(wire_54));
  TC_Switch # (.UUID(64'd4153623403708032652 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_14), .in(wire_69[7:0]), .out(wire_4_8));
  TC_Switch # (.UUID(64'd340002077875967615 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_19), .in(wire_69[7:0]), .out(wire_28_4));
  TC_Or # (.UUID(64'd4530764934882597393 ^ UUID), .BIT_WIDTH(64'd1)) Or_21 (.in0(wire_14), .in1(wire_19), .out(wire_46));
  TC_Or # (.UUID(64'd3471186985449771457 ^ UUID), .BIT_WIDTH(64'd1)) Or_22 (.in0(wire_35), .in1(wire_6), .out(wire_17));
  TC_Ram # (.UUID(64'd4536271034189926213 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_23 (.clk(clk), .rst(rst), .load(wire_46), .save(wire_6), .address({{24{1'b0}}, wire_7 }), .in0({{56{1'b0}}, wire_0 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_69), .out1(), .out2(), .out3());
  TC_Or # (.UUID(64'd1292995358292959653 ^ UUID), .BIT_WIDTH(64'd1)) Or_24 (.in0(wire_13), .in1(wire_39), .out(wire_40));
  TC_Program # (.UUID(64'd4309608288760828634 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_3BCECDE7C4AB12DA.w8.bin"), .ARG_SIG("Program_3BCECDE7C4AB12DA=%s")) Program_25 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_36 }), .out0(wire_27), .out1(wire_10), .out2(wire_5), .out3(wire_38));
  TC_Switch # (.UUID(64'd4415714550226385752 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_26), .in(wire_12), .out(wire_4_5));
  TC_Switch # (.UUID(64'd1189653700547940041 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_23), .in(wire_12), .out(wire_28_3));
  TC_And # (.UUID(64'd155618999696402220 ^ UUID), .BIT_WIDTH(64'd1)) And_28 (.in0(wire_22), .in1(wire_11), .out(wire_25));
  TC_And # (.UUID(64'd541274795936718914 ^ UUID), .BIT_WIDTH(64'd1)) And_29 (.in0(wire_76), .in1(wire_41), .out(wire_21));
  TC_Not # (.UUID(64'd4083299788580941265 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_22), .out(wire_76));
  TC_Or # (.UUID(64'd120137714479852463 ^ UUID), .BIT_WIDTH(64'd1)) Or_31 (.in0(wire_26), .in1(wire_23), .out(wire_41));
  TC_Not # (.UUID(64'd757151366404161751 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_35), .out(wire_33));
  TC_Switch # (.UUID(64'd4421006866021078363 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_33), .in(wire_74), .out(wire_0_0));
  TC_Or # (.UUID(64'd1905578430637404097 ^ UUID), .BIT_WIDTH(64'd1)) Or_34 (.in0(wire_56), .in1(wire_25), .out(wire_2));
  TC_Switch # (.UUID(64'd1874573077821227236 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_56), .in(wire_68), .out(wire_0_1));
  TC_Add # (.UUID(64'd4216442262429427720 ^ UUID), .BIT_WIDTH(64'd8)) Add8_36 (.in0(wire_36), .in1(wire_64), .ci(1'd0), .out(wire_68), .co());
  TC_Constant # (.UUID(64'd3759199946427123610 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_37 (.out(wire_64));
  TC_Splitter8 # (.UUID(64'd4026341976731187117 ^ UUID)) Splitter8_38 (.in(wire_27[7:0]), .out0(), .out1(), .out2(), .out3(wire_50), .out4(wire_43), .out5(wire_62), .out6(wire_32), .out7(wire_66));
  TC_Or # (.UUID(64'd4069589641566867169 ^ UUID), .BIT_WIDTH(64'd1)) Or_39 (.in0(wire_15), .in1(wire_21), .out(wire_31));
  TC_Mux # (.UUID(64'd2849789493388807607 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_40 (.sel(wire_15), .in0(wire_38[7:0]), .in1(wire_12), .out(wire_70));
  TC_And # (.UUID(64'd4463487709450428676 ^ UUID), .BIT_WIDTH(64'd1)) And_41 (.in0(wire_32), .in1(wire_66), .out(wire_63));
  TC_And # (.UUID(64'd4242965850164722796 ^ UUID), .BIT_WIDTH(64'd1)) And_42 (.in0(wire_50), .in1(wire_62), .out(wire_72));
  TC_And # (.UUID(64'd397387688674597742 ^ UUID), .BIT_WIDTH(64'd1)) And_43 (.in0(wire_72), .in1(wire_63), .out(wire_61));
  TC_And # (.UUID(64'd2247596313551031113 ^ UUID), .BIT_WIDTH(64'd1)) And_44 (.in0(wire_48), .in1(wire_61), .out(wire_15));
  TC_And # (.UUID(64'd4041230106421252530 ^ UUID), .BIT_WIDTH(64'd1)) And_45 (.in0(wire_61), .in1(wire_43), .out(wire_56));
  TC_Not # (.UUID(64'd3096427652403559373 ^ UUID), .BIT_WIDTH(64'd1)) Not_46 (.in(wire_43), .out(wire_48));
  TC_Switch # (.UUID(64'd4145945214416329298 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_79), .in(wire_38[7:0]), .out(wire_86));
  TC_Not # (.UUID(64'd2096284966625824862 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_35), .out(wire_79));
  REG # (.UUID(64'd1282751658120047660 ^ UUID)) REG_49 (.clk(clk), .rst(rst), .Load(wire_24), .Input(wire_59), .Save_value(wire_0), .Save(wire_29), .Always_output(wire_7), .Output_1(wire_28_0), .Output_2(wire_4_6));
  REG # (.UUID(64'd3844733500531091050 ^ UUID)) REG_50 (.clk(clk), .rst(rst), .Load(wire_37), .Input(wire_78), .Save_value(wire_0), .Save(wire_49), .Always_output(), .Output_1(wire_28_2), .Output_2(wire_4_4));
  REG # (.UUID(64'd1565800838397152933 ^ UUID)) REG_51 (.clk(clk), .rst(rst), .Load(wire_53), .Input(wire_67), .Save_value(wire_0), .Save(wire_34), .Always_output(), .Output_1(wire_28_5), .Output_2(wire_4_3));
  REG # (.UUID(64'd2505076439785491486 ^ UUID)) REG_52 (.clk(clk), .rst(rst), .Load(wire_84), .Input(wire_55), .Save_value(wire_0), .Save(wire_82), .Always_output(), .Output_1(wire_28_6), .Output_2(wire_4_0));
  REG # (.UUID(64'd120818865867497515 ^ UUID)) REG_53 (.clk(clk), .rst(rst), .Load(wire_30), .Input(wire_81), .Save_value(wire_0), .Save(wire_85), .Always_output(), .Output_1(wire_28_8), .Output_2(wire_4_1));
  ALU # (.UUID(64'd3501525809347837570 ^ UUID)) ALU_54 (.clk(clk), .rst(rst), .Instruction(wire_27[7:0]), .Input_1(wire_58), .Input_2(wire_1), .Output(wire_74));
  DEC # (.UUID(64'd3684352349505994725 ^ UUID)) DEC_55 (.clk(clk), .rst(rst), .Input(wire_27[7:0]), .Output_1(wire_18), .Output_2(wire_16));
  COND # (.UUID(64'd1443519742035116363 ^ UUID)) COND_56 (.clk(clk), .rst(rst), .\4 (wire_52), .\2 (wire_60), .\1 (wire_71), .ARG1(wire_58), ._ARG2(wire_1), .Output(wire_44));
  STACK # (.UUID(64'd957653762625945146 ^ UUID)) STACK_57 (.clk(clk), .rst(rst), .POP(wire_31), .PUSH(wire_2), .VALUE(wire_0), .OUTPUT(wire_12));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  assign wire_0 = wire_0_0|wire_0_1;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  wire [7:0] wire_4_4;
  wire [7:0] wire_4_5;
  wire [7:0] wire_4_6;
  wire [7:0] wire_4_7;
  wire [7:0] wire_4_8;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7|wire_4_8;
  wire [63:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [63:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [63:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_28_0;
  wire [7:0] wire_28_1;
  wire [7:0] wire_28_2;
  wire [7:0] wire_28_3;
  wire [7:0] wire_28_4;
  wire [7:0] wire_28_5;
  wire [7:0] wire_28_6;
  wire [7:0] wire_28_7;
  wire [7:0] wire_28_8;
  assign wire_28 = wire_28_0|wire_28_1|wire_28_2|wire_28_3|wire_28_4|wire_28_5|wire_28_6|wire_28_7|wire_28_8;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [63:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  assign arch_input_enable = wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [7:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [63:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  assign arch_output_enable = wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [7:0] wire_86;
  wire [0:0] wire_87;

endmodule
